* C:\Users\raiha\OneDrive\Desktop\Courses\CSE250\Practice pspice\Schematic1.sch

* Schematics Version 9.1 - Web Update 1
* Sat Nov 20 03:55:31 2021



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic1.net"
.INC "Schematic1.als"


.probe


.END
